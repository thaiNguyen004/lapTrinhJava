�� sr main.sinhVien�1l�% D diemTrungBinhI tuoiL 
maSinhVient Ljava/lang/String;L tenSinhVienq ~ xp@#������   t 001t Nguyênsq ~  @"         t 003t Vinh